module and(
  input a,b,
  output c
);
  and(c,a,b);
endmodule
