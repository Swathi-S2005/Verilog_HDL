module tb;
reg [13*8:1]s;
initial begin
s="hello world";
$display("value of s=%s",s[104:65]);
end
endmodule

