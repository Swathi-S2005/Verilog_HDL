module xorgate(
input a,b,
output y);
xor g1(c,a,b);
endmodule

