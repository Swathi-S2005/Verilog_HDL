module and_gate(
input a,b,
output o);
and g(o,a,b);
endmodule

