module notgate(
input a,en,
output y);
notif1 n1(y,a,en);
endmodule
         
