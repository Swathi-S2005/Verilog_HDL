module notgate(
input a,
output y);
assign y= ~a;
endmodule

