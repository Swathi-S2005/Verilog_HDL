module demux(
input a,s,
output y0,y1);

