module notgate(
input a,en,
output y);
notif0 n1(y,a,en);
endmodule
