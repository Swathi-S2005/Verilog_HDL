module tb_
