module tb_xor;
reg a,b;
wire y;
xorgate uut(
.a(a),
.b(b),
.y(y));
initial begin
$dumpfile("xorgate.vcd");
$dumpvars(0,tb_xor);
$monitor("Time=%0t|a=%b|b=%b|y=%b",$time,a,b,y);
a=0;b=0;#10;
a=0;a=1;#10;
a=1;b=0;#10;
a=1;b=1;#10;
$finish;
end
endmodule

