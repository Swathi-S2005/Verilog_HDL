module notgate(
	input a,
output y);
not g1(y,a);
endmodule

