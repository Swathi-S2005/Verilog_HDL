module int;
integer b;
initial
begin
b= -'d12/3;
end
initial begin
$display("b=%d",b);
end
endmodule
