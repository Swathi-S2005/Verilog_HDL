module nandgate(
input a,b,
output y);
nand g1(y,a,b);
endmodule

